----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.04.2024 22:43:30
-- Design Name: 
-- Module Name: Add_Sub_4bit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Add_Sub_4bit is
    Port ( A : in STD_LOGIC_VECTOR (3 downto 0);
           B : in STD_LOGIC_VECTOR (3 downto 0);
           M : in STD_LOGIC;
           S : out STD_LOGIC_VECTOR (3 downto 0);
           C_out : out STD_LOGIC;
           Overflow : out STD_LOGIC;
           Sign: out STD_LOGIC;
           Zero : out STD_LOGIC );
           
end Add_Sub_4bit;

architecture Behavioral of Add_Sub_4bit is

component FA   
            port (      
            A: in std_logic;     
            B: in std_logic;   
            C_in: in std_logic;  
            S: out std_logic;     
            C_out: out std_logic); 
     end component; 
     
signal FA0_C, FA1_C, FA2_C, FA3_C  : std_logic; 
signal TMP: std_logic_vector(3 downto 0);
signal sum: std_logic_vector(3 downto 0);
signal C_output:  std_logic; 

begin

FA_0 : FA         
    port map (               
        A => A(0),               
        B => TMP(0),             
        C_in => M,        
        S => sum(0),               
        C_out => FA0_C);       
 FA_1 : FA         
    port map (              
        A => A(1),               
        B => TMP(1),             
        C_in => FA0_C,                
        S => sum(1),               
        C_out => FA1_C);    
     
FA_2 : FA         
     port map (               
        A => A(2),               
        B => TMP(2),             
        C_in => FA1_C,                
        S => sum(2),               
        C_out => FA2_C);      
FA_3 : FA         
     port map (               
        A => A(3),               
        B => TMP(3),             
        C_in => FA2_C,                
        S => sum(3),               
        C_out => C_output); 
        
TMP(0)<= M XOR B(0);
TMP(1)<= M XOR B(1);
TMP(2)<= M XOR B(2);
TMP(3)<= M XOR B(3);

C_out<=C_output;
S<=sum; 

Overflow <= FA2_C XOR C_output;
Zero <= (NOT sum(0)) AND (NOT sum(1)) AND (NOT sum(2)) AND (NOT sum(3));
Sign<=sum(3);

end Behavioral;
