----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 13.04.2024 13:03:34
-- Design Name: 
-- Module Name: Mux_2_way_4_bit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Mux_2_way_4_bit is
    Port ( S : in STD_LOGIC;
           A : in STD_LOGIC_VECTOR (3 downto 0);
           B : in STD_LOGIC_VECTOR (3 downto 0);
           Y : out STD_LOGIC_VECTOR (3 downto 0));
end Mux_2_way_4_bit;

architecture Behavioral of Mux_2_way_4_bit is

signal Y0,Y1,Y2,Y3 : STD_LOGIC;

begin

Y0 <= ((A(0) AND (NOT S)) OR (B(0) AND S));
Y1 <= ((A(1) AND (NOT S)) OR (B(1) AND S));
Y2 <= ((A(2) AND (NOT S)) OR (B(2) AND S));
Y3 <= ((A(3) AND (NOT S)) OR (B(3) AND S));
   
Y(0) <= Y0;
Y(1) <= Y1;
Y(2) <= Y2;
Y(3) <= Y3;

end Behavioral;
